//-------------------------------------------------------------------------
//    mb_usb_hdmi_top.sv                                                 --
//    Zuofu Cheng                                                        --
//    2-29-24                                                            --
//                                                                       --
//                                                                       --
//    Spring 2024 Distribution                                           --
//                                                                       --
//    For use with ECE 385 USB + HDMI                                    --
//    University of Illinois ECE Department                              --
//-------------------------------------------------------------------------


module mb_usb_hdmi_top(
    input logic Clk,
    input logic reset_rtl_0,
    
    //USB signals
    input logic [0:0] gpio_usb_int_tri_i,
    output logic gpio_usb_rst_tri_o,
    input logic usb_spi_miso,
    output logic usb_spi_mosi,
    output logic usb_spi_sclk,
    output logic usb_spi_ss,
    
    //UART
    input logic uart_rtl_0_rxd,
    output logic uart_rtl_0_txd,
    
    //HDMI
    output logic hdmi_tmds_clk_n,
    output logic hdmi_tmds_clk_p,
    output logic [2:0]hdmi_tmds_data_n,
    output logic [2:0]hdmi_tmds_data_p,
        
    //HEX displays
    output logic [7:0] hex_segA,
    output logic [3:0] hex_gridA,
    output logic [7:0] hex_segB,
    output logic [3:0] hex_gridB
);
    
    logic [31:0] keycode0_gpio, keycode1_gpio;
    logic clk_25MHz, clk_125MHz, clk_100MHz;
    logic locked;
    logic [9:0] drawX, drawY, ballxsig, ballysig, ballsizesig, knifexsig, knifeysig, knifesizesig;
    logic [9:0] fireballxsig, fireballysig, fireballsizesig;
    logic hsync, vsync, vde;
    logic [3:0] red, green, blue;
    logic reset_ah;

    //World Map
    logic [28:0] info_ground[16], info_ground_0[16], info_ground_1[16];
    logic [28:0] info_fence[16], info_fence_0[16], info_fence_1[16];
    logic [9:0] info_exit[2], info_exit_0[2], info_exit_1[2];
    logic [20:0] info_spince[6], info_spince_0[6], info_spince_1[6];
    logic [20:0] info_monster, info_monster_0, info_monster_1;

    //Logic Block
    logic logic_in_air;
    logic touch_down, touch_up, touch_left, touch_right;
    logic go_up, go_left, go_right;
    logic [9:0] touch_down_position_y, touch_up_position_y, touch_left_position_x, touch_right_position_x;
    logic knife_touch_fence;  
    //win or lose
    logic win_the_game, lose_the_game;

    //state machine
    logic [3:0] game_state;
    logic [1:0] selector_value;

    //monster
    logic monster_exist, fireball_exist;

    assign reset_ah = reset_rtl_0;
    
    
    //Keycode HEX drivers
    hex_driver HexA (
        .clk(Clk),
        .reset(reset_ah),
        .in({keycode0_gpio[31:28], keycode0_gpio[27:24], keycode0_gpio[23:20], keycode0_gpio[19:16]}),
        .hex_seg(hex_segA),
        .hex_grid(hex_gridA)
    );
    
    hex_driver HexB (
        .clk(Clk),
        .reset(reset_ah),
        .in({keycode0_gpio[15:12], keycode0_gpio[11:8], keycode0_gpio[7:4], keycode0_gpio[3:0]}),
        .hex_seg(hex_segB),
        .hex_grid(hex_gridB)
    );
    
    mb_block mb_block_i (
        .clk_100MHz(Clk),
        .gpio_usb_int_tri_i(gpio_usb_int_tri_i),
        .gpio_usb_keycode_0_tri_o(keycode0_gpio),
        .gpio_usb_keycode_1_tri_o(keycode1_gpio),
        .gpio_usb_rst_tri_o(gpio_usb_rst_tri_o),
        .reset_rtl_0(~reset_ah), //Block designs expect active low reset, all other modules are active high
        .uart_rtl_0_rxd(uart_rtl_0_rxd),
        .uart_rtl_0_txd(uart_rtl_0_txd),
        .usb_spi_miso(usb_spi_miso),
        .usb_spi_mosi(usb_spi_mosi),
        .usb_spi_sclk(usb_spi_sclk),
        .usb_spi_ss(usb_spi_ss)
    );
        
    //clock wizard configured with a 1x and 5x clock for HDMI
    clk_wiz_0 clk_wiz (
        .clk_out1(clk_25MHz),
        .clk_out2(clk_125MHz),
        .reset(reset_ah),
        .locked(locked),
        .clk_in1(Clk)
    );
    
    //VGA Sync signal generator
    vga_controller vga (
        .pixel_clk(clk_25MHz),
        .reset(reset_ah),
        .hs(hsync),
        .vs(vsync),
        .active_nblank(vde),
        .drawX(drawX),
        .drawY(drawY)
    );    

    //Real Digital VGA to HDMI converter
    hdmi_tx_0 vga_to_hdmi (
        //Clocking and Reset
        .pix_clk(clk_25MHz),
        .pix_clkx5(clk_125MHz),
        .pix_clk_locked(locked),
        //Reset is active LOW
        .rst(reset_ah),
        //Color and Sync Signals
        .red(red),
        .green(green),
        .blue(blue),
        .hsync(hsync),
        .vsync(vsync),
        .vde(vde),
        
        //aux Data (unused)
        .aux0_din(4'b0),
        .aux1_din(4'b0),
        .aux2_din(4'b0),
        .ade(1'b0),
        
        //Differential outputs
        .TMDS_CLK_P(hdmi_tmds_clk_p),          
        .TMDS_CLK_N(hdmi_tmds_clk_n),          
        .TMDS_DATA_P(hdmi_tmds_data_p),         
        .TMDS_DATA_N(hdmi_tmds_data_n)          
    );

    
    //Ball Module
    ball ball_instance(
        .Reset(reset_ah),
        .frame_clk(vsync),                    //Figure out what this should be so that the ball will move
        .keycode(keycode0_gpio),    //Notice: only one keycode connected to ball by default
        .BallX(ballxsig),
        .BallY(ballysig),
        .BallS(ballsizesig),
        .game_state(game_state),
        .logic_in_air(logic_in_air),
        .touch_down(touch_down),
        .touch_up(touch_up),
        .touch_left(touch_left),
        .touch_right(touch_right),
        .touch_down_position_y(touch_down_position_y),
        .touch_up_position_y(touch_up_position_y),
        .touch_left_position_x(touch_left_position_x),
        .touch_right_position_x(touch_right_position_x),
        .go_up(go_up),
        .go_left(go_left),
        .go_right(go_right)
    );
    
    //Knife Module
    knife knife_instance(
        .Reset(reset_ah),
        .frame_clk(vsync),
        .keycode(keycode0_gpio),
        .BallX(ballxsig),
        .BallY(ballysig),
        .BallS(ballsizesig),
        .go_left(go_left),
        .go_right(go_right),
        .knifeX(knifexsig),
        .knifeY(knifeysig),
        .knifeS(knifesizesig),
        .knife_touch_fence(knife_touch_fence)
    );

    //Color Mapper Module   
    color_mapper color_instance(
        .Clk(clk_25MHz),
        .vde(vde),
        .BallX(ballxsig),
        .BallY(ballysig),
        .DrawX(drawX),
        .DrawY(drawY),
        .Ball_size(ballsizesig),
        .Red(red),
        .Green(green),
        .Blue(blue),
        .info_ground(info_ground),
        .info_fence(info_fence),
        .info_exit(info_exit),
        .info_spince(info_spince),
        .KnifeX(knifexsig),
        .KnifeY(knifeysig),
        .Knife_size(knifesizesig),
        .go_left(go_left),
        .go_right(go_right),
        .game_state(game_state),
        .fireballX(fireballxsig),
        .fireballY(fireballysig),
        .fireballS(fireballsizesig),
        .fireball_exist(fireball_exist),
        .monster_exist(monster_exist),
        .info_monster(info_monster)
    );

    world_map world_map_instance(
        .Reset(reset_ah),
        .Clk(vsync),
        .info_ground(info_ground_1),
        .info_fence(info_fence_1),
        .info_exit(info_exit_1),
        .info_spince(info_spince_1),
        .BallX(ballxsig),
        .BallY(ballysig),
        .info_monster(info_monster_1),
        .monster_exist(monster_exist)
    );

    world_map_0 world_map_0_instance(
        .Reset(reset_ah),
        .Clk(vsync),
        .info_ground(info_ground_0),
        .info_fence(info_fence_0),
        .info_exit(info_exit_0),
        .info_spince(info_spince_0),
        .BallX(ballxsig),
        .BallY(ballysig),
        .info_monster(info_monster_0),
        .monster_exist(monster_exist)
    );

    logic_block logic_block_instance(
        .pixel_clk(vsync),
        .reset(reset_ah),
        .BallX(ballxsig),
        .BallY(ballysig),
        .BallS(ballsizesig),
        .KnifeX(knifexsig),
        .KnifeY(knifeysig),
        .KnifeS(knifesizesig),
        .logic_in_air(logic_in_air),
        .info_ground(info_ground),
        .info_fence(info_fence),
        .info_exit(info_exit),
        .info_spince(info_spince),
        .touch_down(touch_down),
        .touch_up(touch_up),
        .touch_left(touch_left),
        .touch_right(touch_right),
        .knife_touch_fence(knife_touch_fence),
        .touch_down_position_y(touch_down_position_y),
        .touch_up_position_y(touch_up_position_y),
        .touch_left_position_x(touch_left_position_x),
        .touch_right_position_x(touch_right_position_x),
        .go_up(go_up),
        .go_left(go_left),
        .go_right(go_right),
        .win_the_game(win_the_game),
        .lose_the_game(lose_the_game),
        .fireballX(fireballxsig),
        .fireballY(fireballysig),
        .fireballS(fireballsizesig)
    );

    state_machine state_machine_instance(
        .reset(reset_ah),
        .pixel_clk(vsync),
        .game_state(game_state),
        .keycode(keycode0_gpio),
        .win_the_game(win_the_game),
        .lose_the_game(lose_the_game),
        .selector_value(selector_value)
    );

    world_selector world_selector_instance(
        .Reset(reset_ah),
        .Clk(vsync),
        .selector_value(selector_value),
        
        .info_ground_0(info_ground_0),
        .info_fence_0(info_fence_0),
        .info_exit_0(info_exit_0),
        .info_spince_0(info_spince_0),
        .info_monster_0(info_monster_0),
        
        .info_ground_1(info_ground_1),
        .info_fence_1(info_fence_1),
        .info_exit_1(info_exit_1),
        .info_spince_1(info_spince_1),
        .info_monster_1(info_monster_1),
        
        .info_ground(info_ground),
        .info_fence(info_fence),
        .info_exit(info_exit),
        .info_spince(info_spince),
        .info_monster(info_monster)
    );

    monster monster_instance(
        .Reset(reset_ah),
        .frame_clk(vsync),
        .BallX(ballxsig),
        .BallY(ballysig),
        .BallS(ballsizesig),
        .info_monster(info_monster),
        .game_state(game_state),
        .fireballX(fireballxsig),
        .fireballY(fireballysig),
        .fireballS(fireballsizesig),
        .fireball_exist(fireball_exist),
        .knifeX(knifexsig),
        .knifeY(knifeysig),
        .monster_exist(monster_exist)
    );

 
endmodule
