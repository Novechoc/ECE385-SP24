/*
 * ECE385-HelperTools/PNG-To-Txt
 * Author: Rishi Thakkar
 *
 */

module  frameRAM
(
		input [18:0]read_address,
		input Clk,

		output logic [3:0] data_Out
);

// mem has width of 3 bits and a total of 400 addresses
logic [3:0] mem [0:30719];

initial
begin
	 $readmemh("ram_file/123.txt", mem);
end


always_comb begin
	data_Out<= mem[read_address];
end

endmodule
